`ifndef DICE_DEFINE_VH
`define DICE_DEFINE_VH

`include "dice_config.vh"

`endif // DICE_DEFINE_VH
