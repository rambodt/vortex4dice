// tcu_pkg.sv
package tcu_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;

  //------------------------------------------
  // Transaction Items
  //------------------------------------------
  `include "tcu_seq_item.svh"
  `include "tcu_out_item.svh"

  //------------------------------------------
  // Agent Components
  //------------------------------------------
  `include "tcu_driver.svh"
  `include "tcu_monitor.svh"
  `include "tcu_sequencer.svh"
  `include "tcu_agent.svh"

  //------------------------------------------
  // Sequences
  //------------------------------------------
  `include "tcu_random_seq.svh"

  //------------------------------------------
  // Environment Components
  //------------------------------------------
  `include "tcu_scoreboard.svh"
  `include "tcu_env.svh"

  //------------------------------------------
  // Tests
  //------------------------------------------
  `include "tcu_base_test.svh"

endpackage